library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity FIFO8x9 is
   port(
      clk, rst:		in std_logic;
      RdPtrClr, WrPtrClr:	in std_logic;    
      RdInc, WrInc:	in std_logic;
      DataIn:	 in std_logic_vector(8 downto 0);
      DataOut: out std_logic_vector(8 downto 0);
      rden, wren: in std_logic
	);
end entity FIFO8x9;

architecture RTL of FIFO8x9 is
	--signal declarations
	type fifo_array is array(7 downto 0) of std_logic_vector(8 downto 0);  -- makes use of VHDL’s enumerated type
	signal fifo:  fifo_array;
	signal wrptr, rdptr: unsigned(2 downto 0);
	signal en: std_logic_vector(7 downto 0);
	signal dmuxout: std_logic_vector(8 downto 0);
begin
process (clk,rst) begin
	if rst = '1' then 
		for i in 7 downto 0 loop
			fifo(i) <= "000000000";
			wrptr <= "000";
			rdptr <= "000";
		end loop;
	elsif rising_edge(clk) then
			if rden = '1' then 
				DataOut <= fifo(to_integer(unsigned(rdptr))) ;
			else 
				DataOut <= "ZZZZZZZZZ";
			end if;
			if wren = '1' then
				fifo(to_integer(unsigned(wrptr))) <= DataIn;
                        else
				fifo(to_integer(unsigned(wrptr))) <= fifo(to_integer(unsigned(wrptr)));
                        end if;
	if WrPtrClr = '0' then
		wrptr <= "000";
	elsif RdInc = '1' then
		wrptr <= wrptr +1;
	end if;
	if WrPtrClr = '0' then
		wrptr <= "000";
	elsif WrInc = '1' then
		wrptr <= wrptr +1;
	end if;
			
	end if;
 



end process;
end RTL;
